// ----  Probes  ----
`define PROBE_ADDR       probe_addr
`define PROBE_DATA_IN    probe_data_in
`define PROBE_DATA_OUT   mem_data_out
`define PROBE_READ_EN    probe_read_en
`define PROBE_WRITE_EN   probe_write_en

`define PROBE_F_PC       u_fetch.pc_o
`define PROBE_F_INSN     u_fetch.insn_o
// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd1
// ----  Top module  ----

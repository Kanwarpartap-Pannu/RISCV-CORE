`define PROBE_ADDR      mem_addr
`define PROBE_DATA_IN   mem_data_in
`define PROBE_DATA_OUT  mem_data_out
`define PROBE_READ_EN   mem_read_en
`define PROBE_WRITE_EN  mem_write_en

`define PROBE_F_PC      f_pc
`define PROBE_F_INSN    f_insn

// ----  Top module  ----
`define TOP_MODULE  pd1
// ----  Top module  ----